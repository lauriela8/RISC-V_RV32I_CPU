`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:2**8-1];

    initial begin
        //$readmemh("code.mem", rom);

        // R-Type  funct7(7) | rs2(5) | rs1(5) | funct3(3) | rd(5) | opcode(7)
        rom[0]  = 32'b0000000_00010_00001_000_00100_0110011; // add   x4,  x1, x2
        rom[1]  = 32'b0100000_00010_00001_000_00101_0110011; // sub   x5,  x1, x2
        rom[2]  = 32'b0000000_00010_00001_001_00110_0110011; // sll   x6,  x1, x2
        rom[3]  = 32'b0000000_00010_00001_010_00111_0110011; // slt   x7,  x1, x2
        rom[4]  = 32'b0000000_00010_00001_011_01000_0110011; // sltu  x8,  x1, x2
        rom[5]  = 32'b0000000_00010_00001_100_01001_0110011; // xor   x9,  x1, x2
        rom[6] = 32'b0000000_00010_00001_101_01010_0110011; // srl   x10, x1, x2
        rom[7] = 32'b0100000_00010_00001_101_01011_0110011; // sra   x11, x1, x2
        rom[8] = 32'b0000000_00010_00001_110_01100_0110011; // or    x12, x1, x2
        rom[9] = 32'b0000000_00010_00001_111_01101_0110011; // and   x13, x1, x2

        // I-Type  imm[11:0](12) | rs1(5) | funct3(3) | rd(5) | opcode(7)
        rom[10] = 32'b000000000100_00001_000_01110_0010011;  // addi  x14, x1, 4
        rom[11] = 32'b000000000100_00001_010_01111_0010011;  // slti  x15, x1, 4
        rom[12] = 32'b000000000100_00001_011_10000_0010011;  // sltiu x16, x1, 4
        rom[13] = 32'b000000000100_00001_100_10001_0010011;  // xori  x17, x1, 4
        rom[14] = 32'b000000000100_00001_110_10010_0010011;  // ori   x18, x1, 4
        rom[15] = 32'b000000000100_00001_111_10011_0010011;  // andi  x19, x1, 4
        rom[16] = 32'b0000000_00010_00001_001_10100_0010011; // slli  x20, x1, x2
        rom[17] = 32'b0000000_00010_00001_101_10101_0010011; // srli  x21, x1, x2
        rom[18] = 32'b0100000_00010_00001_101_10110_0010011; // srai  x22, x1, x2

        // S-Type  imm[11:5](7) | rs2(5) | rs1(5) | funct3(3) | imm[4:0](5) | opcode(7)
        rom[19] = 32'b0000000_00100_00001_010_00000_0100011;  // sw x4, 0(x1)
        rom[20] = 32'b0000000_00101_00001_000_00100_0100011;  // sb x5, 4(x1)
        rom[21] = 32'b0000000_00110_00001_001_01000_0100011;  // sh x6, 8(x1)

        // L-Type  imm[11:0](12) | rs1(5) | funct3(3) | rd(5) | opcode(7)
        rom[22] = 32'b000000000000_00001_000_10111_0000011;  // lb  x23, 0(x1)
        rom[23] = 32'b000000000100_00001_001_11000_0000011;  // lh  x24, 4(x1)
        rom[24] = 32'b000000001000_00001_010_11001_0000011;  // lw  x25, 8(x1)
        rom[25] = 32'b000000000100_00001_100_11010_0000011;  // lbu x26, 4(x1)
        rom[26] = 32'b000000001000_00001_101_11011_0000011;  // lhu x27, 8(x1)

        rom[27] = 32'b0000000_00001_00001_000_00100_1100011;  // beq   x1, x1, +4
        rom[28] = 32'b0000000_00010_00001_001_00100_1100011;  // bne   x1, x2, +4
        rom[29] = 32'b0000000_00001_00010_100_00100_1100011;  // blt   x1, x2, +4
        rom[30] = 32'b0000000_00001_00010_101_00100_1100011;  // bge   x1, x2, +4
        rom[31] = 32'b0000000_00001_00010_110_00100_1100011; // bltu  x1, x2, +4
        rom[32] = 32'b0000000_00001_00010_111_00100_1100011; // bgeu  x1, x2, +4

        // U-Type  imm[31:12](20) | rd(5) | opcode(7)
        rom[33] = 32'b00000000000000000001_11100_0110111;  // lui   x28, 1
        rom[34] = 32'b00000000000000000001_11101_0010111;  // auipc x29, 1

        rom[35] = 32'b0_0000000001_0_00000000_11110_1101111;  // jal  x30, +4
        rom[36] = 32'b000000000100_00001_000_11111_1100111;  // jalr x31, 4(x1)

        // J-Type  imm[20|10:1|11|19:12](20) | rd(5) | opcode(7)
        //rom[33] = 32'b0_0000000100_0_00000000_11110_1101111; // jal x30, 8           

        // J-Type (JALR)  imm[11:0](12) | rs1(5) | funct3(3) | rd(5) | opcode(7)
        //rom[35] = 32'b000010001100_00100_000_11111_1100111;  // jalr x31, x4, 140

    end

    assign data = rom[addr[31:2]];
endmodule
