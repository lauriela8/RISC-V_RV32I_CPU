`timescale 1ns / 1ps

module MCU (
    input logic clk,
    input logic rst
);
    logic [31:0] instrCode;
    logic [31:0] instrMemAddr;
    logic        busWe;
    logic [31:0] busAddr;
    logic [31:0] busWData;
    logic [31:0] busRData;
    logic [ 2:0] busFunc3;

    ROM U_ROM (
        .addr(instrMemAddr),
        .data(instrCode)
    );

    CPU_RV32I U_RV32I (.*);

    RAM U_RAM (
        .clk  (clk),
        .we   (busWe),
        .func3(busFunc3),
        .addr (busAddr),
        .wData(busWData),
        .rData(busRData)
    );
endmodule
